module seven_segment(
	input [7:0] digital_signal,
	output [6:0] segments,
	output [2:0] digit_select
	);
	
	
	
endmodule